LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY aula10_exercicio1 IS
	PORT(SW   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		  HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6));	
END ENTITY;

ARCHITECTURE dec_bcd OF aula10_exercicio1 IS
BEGIN
	PROCESS(SW)
	BEGIN
		CASE SW IS
			WHEN "0000" => HEX0 <= "0000001"; --0
			WHEN "0001" => HEX0 <= "1001111"; --1
			WHEN "0010" => HEX0 <= "0010010"; --2
			WHEN "0011" => HEX0 <= "0000110"; --3
			WHEN "0100" => HEX0 <= "1001100"; --4
			WHEN "0101" => HEX0 <= "0100100"; --5
			WHEN "0110" => HEX0 <= "0100000"; --6
			WHEN "0111" => HEX0 <= "0001111"; --7
			WHEN "1000" => HEX0 <= "0000000"; --8
			WHEN "1001" => HEX0 <= "0000100"; --9
			WHEN OTHERS => HEX0 <= "0110000"; --E
		END CASE;
	END PROCESS;
END ARCHITECTURE;
