LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula11_exercicio1 IS
	GENERIC (N : INTEGER := 4);
	PORT(Se  : IN  	STD_LOGIC;
		  CLK : IN  	STD_LOGIC;
		  Q 	: BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE logic OF Aula11_exercicio1 IS
BEGIN
	PROCESS(CLK)
	BEGIN
		FOR i IN 0 TO N-2 LOOP
			IF(CLK'EVENT AND CLK = '1') THEN
				Q(i) <= Q(i + 1);
			END IF;
			Q(N-1) <= Se;
		END LOOP;
	END PROCESS;
	
END;