LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY VHDL_Exemplo2 IS
	PORT (S1 : IN std_logic;
			S2 : IN std_logic;
			A	: IN std_logic;
			B  : IN std_logic;
			C  : IN std_logic;
			D  : IN std_logic;
	  SAIDA : OUT std_logic);
END VHDL_Exemplo2;

ARCHITECTURE logica OF VHDL_Exemplo2 IS 
BEGIN
	SAIDA <= (A AND (NOT S1) AND (NOT S2)) OR
				(B AND (NOT S1) AND S2) OR
				(C AND S1 AND (NOT S2)) OR
				(D AND S1 AND S2);
END logica;
			