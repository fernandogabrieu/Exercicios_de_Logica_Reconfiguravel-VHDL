LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula11_exercicio4 IS
	PORT(A : IN  INTEGER RANGE 0 TO 7;
		  Z :	OUT STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000");
END ENTITY;

ARCHITECTURE logic OF Aula11_exercicio4 IS
BEGIN
	PROCESS
	BEGIN
		WAIT UNTIL A = 2;
		Z <= "1111";
	END PROCESS;
END ARCHITECTURE;