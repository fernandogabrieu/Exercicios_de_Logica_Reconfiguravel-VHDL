LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula11_exercicio3 IS
	PORT(A :  IN INTEGER RANGE 0 TO 7;
		  Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE logic OF Aula11_exercicio3 IS
BEGIN
	PROCESS(A)
		VARIABLE I : INTEGER RANGE 0 TO 4;
	BEGIN
		Z <= "0000";
		I := 0;
		WHILE (I <= 3) LOOP
			IF (A = I) THEN
				Z(I) <= '1';
			END IF;
			I := I + 1;
		END LOOP;
	END PROCESS;
END;