LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY aula10_exercicio4 IS
	PORT(KEY  : STD_LOGIC_VECTOR(0 DOWNTO 0);
		  LEDR : STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE seq_leds OF aula10_exercicio4 IS
BEGIN
	PROCESS(KEY)
	BEGIN
		IF(KEY(0)'EVENT AND KEY(0) = '1') THEN
			CASE KEY IS
				WHEN 
			
		END IF;
	END PROCESS;
END;