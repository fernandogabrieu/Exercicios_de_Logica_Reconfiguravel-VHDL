LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Aula12_Exercicio4 IS
	PORT();
END ENTITY;

ARCHITECTURE logic OF Aula12_Exercicio4 IS
BEGIN└
	PROCESS(clk)
	BEGIN
	END PROCESS;
END;